** Profile: "SCHEMATIC1-Lab5Sim"  [ E:\Circuits-I\Lab5\Lab5-PSpiceFiles\SCHEMATIC1\Lab5Sim.sim ] 

** Creating circuit file "Lab5Sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\cel8473\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1m 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
